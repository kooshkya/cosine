module CUD (input start, clk, rst, input [15:0] v, angle, output done, output [15:0] distance);
    
endmodule